module valve

struct ICvar {}
