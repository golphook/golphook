module valve
//
// import utils
//
// struct ISurface {}
//
// type P_lock_cursor = fn ()
// type P_unlock_cursor = fn ()
//
// pub fn (mut i ISurface) lock_cursor() {
// 	o_fn_add := utils.get_virtual(i, 66)
//
// 	o_fn := &P_lock_cursor(o_fn_add)
// 	o_fn()
// }
//
// pub fn (mut i ISurface) unlock_cursor() {
// 	o_fn_add := utils.get_virtual(i, 67)
//
// 	o_fn := &P_unlock_cursor(o_fn_add)
// 	//load_this(i)
// 	o_fn()
// }
