module valve

struct ICvar {

}
