module valve
//
// import utils
//
// struct UIEngine {}
//
// type P_access_engine = fn() &UIEngine
//
// pub fn (mut u UIEngine) access_engine() &UIEngine {
// 	o_fn_add := utils.get_virtual(i, 11)
//
// 	o_fn := &P_access_engine(o_fn_add)
// 	C.load_this(u)
//
// 	rs := o_fn()
// 	return rs
// }
//
// struct IPanoramaUIEngine {}
//
// type P_access_engine = fn() &UIEngine
//
// pub fn (mut i IPanoramaUIEngine) access_engine() &UIEngine {
// 	o_fn_add := utils.get_virtual(i, 11)
//
// 	o_fn := &P_access_engine(o_fn_add)
// 	C.load_this(i)
//
// 	rs := o_fn()
// 	return rs
// }
