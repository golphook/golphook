module valve

struct ICvar {
}
