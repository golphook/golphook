module utils

pub struct Color {
	r u8
	g u8
	b u8
	a u8
}
